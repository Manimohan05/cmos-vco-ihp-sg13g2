* NGSPICE file created from vco.ext - technology: ihp-sg13g2

.subckt vco VPWR VGND vctl Vout
X0 a_542_269# a_745_n2395# a_684_n1958# VGND sg13_lv_nmos ad=0.11p pd=0.94u as=0.17p ps=1.68u w=0.5u l=0.13u
X1 a_7398_n1956# vctl VGND VGND sg13_lv_nmos ad=65.99999f pd=0.74u as=0.102p ps=1.28u w=0.3u l=0.13u
X2 a_4776_351# a_3434_351# a_4909_n217# VGND sg13_lv_nmos ad=0.11p pd=0.94u as=0.17p ps=1.68u w=0.5u l=0.13u
X3 a_4909_n217# vctl VGND VGND sg13_lv_nmos ad=65.99999f pd=0.74u as=0.102p ps=1.28u w=0.3u l=0.13u
X4 a_4771_n2395# a_6113_n2395# a_6051_n2525# VPWR sg13_lv_pmos ad=0.1106p pd=0.945u as=0.11p ps=0.94u w=0.5u l=0.13u
X5 a_2026_n1958# vctl VGND VGND sg13_lv_nmos ad=65.99999f pd=0.74u as=0.102p ps=1.28u w=0.3u l=0.13u
X6 a_6024_351# a_4776_351# Vout VPWR sg13_lv_pmos ad=0.17p pd=1.68u as=0.11p ps=0.94u w=0.5u l=0.13u
X7 a_4909_n217# a_3434_351# a_4776_351# VGND sg13_lv_nmos ad=0.17p pd=1.68u as=0.11p ps=0.94u w=0.5u l=0.13u
X8 a_6113_n2395# Vout a_7397_n2523# VPWR sg13_lv_pmos ad=0.1106p pd=0.945u as=0.11p ps=0.94u w=0.5u l=0.13u
X9 a_656_351# a_542_269# a_750_351# VPWR sg13_lv_pmos ad=0.17p pd=1.68u as=0.11p ps=0.94u w=0.5u l=0.13u
X10 a_7397_n2523# a_620_930# VPWR VPWR sg13_lv_pmos ad=59f pd=0.74u as=0.104p ps=1.34u w=0.2u l=0.13u
X11 VGND vctl a_4909_n217# VGND sg13_lv_nmos ad=0.102p pd=1.28u as=65.99999f ps=0.74u w=0.3u l=0.13u
X12 a_3434_351# VGND cap_cmim l=6.99u w=6.99u
X13 VPWR a_620_930# a_3367_n2525# VPWR sg13_lv_pmos ad=59f pd=0.74u as=59f ps=0.74u w=0.2u l=0.13u
X14 a_3340_351# a_620_930# VPWR VPWR sg13_lv_pmos ad=59.75f pd=0.745u as=0.104p ps=1.34u w=0.2u l=0.13u
X15 a_2092_351# a_750_351# a_1998_351# VPWR sg13_lv_pmos ad=0.11p pd=0.94u as=0.11p ps=0.94u w=0.5u l=0.13u
X16 a_6051_n2525# a_620_930# VPWR VPWR sg13_lv_pmos ad=59f pd=0.74u as=0.104p ps=1.34u w=0.2u l=0.13u
X17 VPWR a_620_930# a_3367_n2525# VPWR sg13_lv_pmos ad=0.104p pd=1.34u as=59.75f ps=0.745u w=0.2u l=0.13u
X18 a_684_n1958# vctl VGND VGND sg13_lv_nmos ad=65.99999f pd=0.74u as=0.102p ps=1.28u w=0.3u l=0.13u
X19 VPWR a_620_930# a_4682_351# VPWR sg13_lv_pmos ad=0.104p pd=1.34u as=59f ps=0.74u w=0.2u l=0.13u
X20 a_683_n2525# a_620_930# VPWR VPWR sg13_lv_pmos ad=59.75f pd=0.745u as=59f ps=0.74u w=0.2u l=0.13u
X21 a_6052_n1958# a_6113_n2395# a_4771_n2395# VGND sg13_lv_nmos ad=0.17p pd=1.68u as=0.11p ps=0.94u w=0.5u l=0.13u
X22 a_2092_351# a_750_351# a_1998_351# VPWR sg13_lv_pmos ad=0.1106p pd=0.945u as=0.17p ps=1.68u w=0.5u l=0.13u
X23 a_7398_n1956# Vout a_6113_n2395# VGND sg13_lv_nmos ad=0.17p pd=1.68u as=0.11p ps=0.94u w=0.5u l=0.13u
X24 VPWR a_620_930# a_3340_351# VPWR sg13_lv_pmos ad=59f pd=0.74u as=59.75f ps=0.745u w=0.2u l=0.13u
X25 a_7397_n2523# Vout a_6113_n2395# VPWR sg13_lv_pmos ad=0.17p pd=1.68u as=0.1106p ps=0.945u w=0.5u l=0.13u
X26 a_2025_n2525# a_2087_n2395# a_745_n2395# VPWR sg13_lv_pmos ad=0.11p pd=0.94u as=0.11p ps=0.94u w=0.5u l=0.13u
X27 VPWR a_620_930# a_4709_n2525# VPWR sg13_lv_pmos ad=59f pd=0.74u as=59f ps=0.74u w=0.2u l=0.13u
X28 a_4709_n2525# a_4771_n2395# a_3429_n2395# VPWR sg13_lv_pmos ad=0.11p pd=0.94u as=0.11p ps=0.94u w=0.5u l=0.13u
X29 VPWR a_620_930# a_2025_n2525# VPWR sg13_lv_pmos ad=0.104p pd=1.34u as=59.75f ps=0.745u w=0.2u l=0.13u
X30 a_2025_n2525# a_2087_n2395# a_745_n2395# VPWR sg13_lv_pmos ad=0.17p pd=1.68u as=0.1106p ps=0.945u w=0.5u l=0.13u
X31 VGND vctl a_6052_n1958# VGND sg13_lv_nmos ad=0.102p pd=1.28u as=65.99999f ps=0.74u w=0.3u l=0.13u
X32 VGND vctl a_7398_n1956# VGND sg13_lv_nmos ad=0.102p pd=1.28u as=65.99999f ps=0.74u w=0.3u l=0.13u
X33 a_6251_n217# a_4776_351# Vout VGND sg13_lv_nmos ad=0.17p pd=1.68u as=0.11p ps=0.94u w=0.5u l=0.13u
X34 VPWR a_620_930# a_7397_n2523# VPWR sg13_lv_pmos ad=59f pd=0.74u as=59f ps=0.74u w=0.2u l=0.13u
X35 VGND vctl a_6251_n217# VGND sg13_lv_nmos ad=0.102p pd=1.28u as=65.99999f ps=0.74u w=0.3u l=0.13u
X36 a_883_n217# a_542_269# a_750_351# VGND sg13_lv_nmos ad=0.17p pd=1.68u as=0.11p ps=0.94u w=0.5u l=0.13u
X37 VGND vctl a_883_n217# VGND sg13_lv_nmos ad=0.102p pd=1.28u as=65.99999f ps=0.74u w=0.3u l=0.13u
X38 VPWR a_620_930# a_3340_351# VPWR sg13_lv_pmos ad=0.104p pd=1.34u as=59f ps=0.74u w=0.2u l=0.13u
X39 a_2092_351# a_750_351# a_2225_n217# VGND sg13_lv_nmos ad=0.11p pd=0.94u as=0.17p ps=1.68u w=0.5u l=0.13u
X40 a_2225_n217# vctl VGND VGND sg13_lv_nmos ad=65.99999f pd=0.74u as=0.102p ps=1.28u w=0.3u l=0.13u
X41 a_3367_n2525# a_3429_n2395# a_2087_n2395# VPWR sg13_lv_pmos ad=0.11p pd=0.94u as=0.11p ps=0.94u w=0.5u l=0.13u
X42 a_4682_351# a_620_930# VPWR VPWR sg13_lv_pmos ad=59f pd=0.74u as=59f ps=0.74u w=0.2u l=0.13u
X43 a_4771_n2395# a_6113_n2395# a_6051_n2525# VPWR sg13_lv_pmos ad=0.11p pd=0.94u as=0.17p ps=1.68u w=0.5u l=0.13u
X44 a_3367_n2525# a_3429_n2395# a_2087_n2395# VPWR sg13_lv_pmos ad=0.17p pd=1.68u as=0.1106p ps=0.945u w=0.5u l=0.13u
X45 a_6024_351# a_620_930# VPWR VPWR sg13_lv_pmos ad=59.75f pd=0.745u as=0.104p ps=1.34u w=0.2u l=0.13u
X46 a_6113_n2395# Vout a_7397_n2523# VPWR sg13_lv_pmos ad=0.11p pd=0.94u as=0.17p ps=1.68u w=0.5u l=0.13u
X47 a_542_269# a_745_n2395# a_683_n2525# VPWR sg13_lv_pmos ad=0.1106p pd=0.945u as=0.11p ps=0.94u w=0.5u l=0.13u
X48 a_3340_351# a_2092_351# a_3434_351# VPWR sg13_lv_pmos ad=0.11p pd=0.94u as=0.1106p ps=0.945u w=0.5u l=0.13u
X49 a_2025_n2525# a_620_930# VPWR VPWR sg13_lv_pmos ad=59f pd=0.74u as=0.104p ps=1.34u w=0.2u l=0.13u
X50 a_745_n2395# a_2087_n2395# a_2025_n2525# VPWR sg13_lv_pmos ad=0.11p pd=0.94u as=0.17p ps=1.68u w=0.5u l=0.13u
X51 a_1998_351# a_620_930# VPWR VPWR sg13_lv_pmos ad=59f pd=0.74u as=59f ps=0.74u w=0.2u l=0.13u
X52 a_542_269# VGND cap_cmim l=6.99u w=6.99u
X53 a_2025_n2525# a_620_930# VPWR VPWR sg13_lv_pmos ad=59.75f pd=0.745u as=59f ps=0.74u w=0.2u l=0.13u
X54 a_656_351# a_620_930# VPWR VPWR sg13_lv_pmos ad=59.75f pd=0.745u as=0.104p ps=1.34u w=0.2u l=0.13u
X55 a_745_n2395# a_2087_n2395# a_2025_n2525# VPWR sg13_lv_pmos ad=0.1106p pd=0.945u as=0.11p ps=0.94u w=0.5u l=0.13u
X56 a_683_n2525# a_620_930# VPWR VPWR sg13_lv_pmos ad=59f pd=0.74u as=0.104p ps=1.34u w=0.2u l=0.13u
X57 a_620_930# vctl VGND VGND sg13_lv_nmos ad=65.99999f pd=0.74u as=0.102p ps=1.28u w=0.3u l=0.13u
X58 a_2087_n2395# a_3429_n2395# a_3368_n1958# VGND sg13_lv_nmos ad=0.11p pd=0.94u as=0.17p ps=1.68u w=0.5u l=0.13u
X59 a_542_269# a_745_n2395# a_683_n2525# VPWR sg13_lv_pmos ad=0.11p pd=0.94u as=0.17p ps=1.68u w=0.5u l=0.13u
X60 VPWR a_620_930# a_4709_n2525# VPWR sg13_lv_pmos ad=0.104p pd=1.34u as=59.75f ps=0.745u w=0.2u l=0.13u
X61 VPWR a_620_930# a_6024_351# VPWR sg13_lv_pmos ad=59f pd=0.74u as=59.75f ps=0.745u w=0.2u l=0.13u
X62 a_684_n1958# a_745_n2395# a_542_269# VGND sg13_lv_nmos ad=0.17p pd=1.68u as=0.11p ps=0.94u w=0.5u l=0.13u
X63 a_1998_351# a_750_351# a_2092_351# VPWR sg13_lv_pmos ad=0.17p pd=1.68u as=0.11p ps=0.94u w=0.5u l=0.13u
X64 VPWR a_620_930# a_656_351# VPWR sg13_lv_pmos ad=59f pd=0.74u as=59.75f ps=0.745u w=0.2u l=0.13u
X65 a_2225_n217# a_750_351# a_2092_351# VGND sg13_lv_nmos ad=0.17p pd=1.68u as=0.11p ps=0.94u w=0.5u l=0.13u
X66 VPWR a_620_930# a_620_930# VPWR sg13_lv_pmos ad=59f pd=0.74u as=59f ps=0.74u w=0.2u l=0.13u
X67 a_3368_n1958# vctl VGND VGND sg13_lv_nmos ad=65.99999f pd=0.74u as=0.102p ps=1.28u w=0.3u l=0.13u
X68 VGND vctl a_2225_n217# VGND sg13_lv_nmos ad=0.102p pd=1.28u as=65.99999f ps=0.74u w=0.3u l=0.13u
X69 a_3429_n2395# VGND cap_cmim l=6.99u w=6.99u
X70 a_3434_351# a_2092_351# a_3340_351# VPWR sg13_lv_pmos ad=0.11p pd=0.94u as=0.11p ps=0.94u w=0.5u l=0.13u
X71 a_3367_n2525# a_620_930# VPWR VPWR sg13_lv_pmos ad=59.75f pd=0.745u as=59f ps=0.74u w=0.2u l=0.13u
X72 a_4682_351# a_620_930# VPWR VPWR sg13_lv_pmos ad=59.75f pd=0.745u as=0.104p ps=1.34u w=0.2u l=0.13u
X73 a_3434_351# a_2092_351# a_3567_n217# VGND sg13_lv_nmos ad=0.11p pd=0.94u as=0.17p ps=1.68u w=0.5u l=0.13u
X74 a_620_930# a_620_930# VPWR VPWR sg13_lv_pmos ad=59f pd=0.74u as=0.104p ps=1.34u w=0.2u l=0.13u
X75 a_2087_n2395# a_3429_n2395# a_3367_n2525# VPWR sg13_lv_pmos ad=0.1106p pd=0.945u as=0.11p ps=0.94u w=0.5u l=0.13u
X76 a_3567_n217# vctl VGND VGND sg13_lv_nmos ad=65.99999f pd=0.74u as=0.102p ps=1.28u w=0.3u l=0.13u
X77 VPWR a_620_930# a_6051_n2525# VPWR sg13_lv_pmos ad=59f pd=0.74u as=59f ps=0.74u w=0.2u l=0.13u
X78 a_3429_n2395# a_4771_n2395# a_4710_n1958# VGND sg13_lv_nmos ad=0.11p pd=0.94u as=0.17p ps=1.68u w=0.5u l=0.13u
X79 VGND vctl a_684_n1958# VGND sg13_lv_nmos ad=0.102p pd=1.28u as=65.99999f ps=0.74u w=0.3u l=0.13u
X80 a_4682_351# a_3434_351# a_4776_351# VPWR sg13_lv_pmos ad=0.11p pd=0.94u as=0.1106p ps=0.945u w=0.5u l=0.13u
X81 a_4771_n2395# VGND cap_cmim l=6.99u w=6.99u
X82 a_6051_n2525# a_6113_n2395# a_4771_n2395# VPWR sg13_lv_pmos ad=0.11p pd=0.94u as=0.11p ps=0.94u w=0.5u l=0.13u
X83 Vout a_4776_351# a_6251_n217# VGND sg13_lv_nmos ad=0.11p pd=0.94u as=0.17p ps=1.68u w=0.5u l=0.13u
X84 a_6251_n217# vctl VGND VGND sg13_lv_nmos ad=65.99999f pd=0.74u as=0.102p ps=1.28u w=0.3u l=0.13u
X85 VPWR a_620_930# a_6024_351# VPWR sg13_lv_pmos ad=0.104p pd=1.34u as=59f ps=0.74u w=0.2u l=0.13u
X86 VPWR a_620_930# a_6051_n2525# VPWR sg13_lv_pmos ad=0.104p pd=1.34u as=59.75f ps=0.745u w=0.2u l=0.13u
X87 a_6051_n2525# a_6113_n2395# a_4771_n2395# VPWR sg13_lv_pmos ad=0.17p pd=1.68u as=0.1106p ps=0.945u w=0.5u l=0.13u
X88 a_3434_351# a_2092_351# a_3340_351# VPWR sg13_lv_pmos ad=0.1106p pd=0.945u as=0.17p ps=1.68u w=0.5u l=0.13u
X89 a_4682_351# a_3434_351# a_4776_351# VPWR sg13_lv_pmos ad=0.17p pd=1.68u as=0.11p ps=0.94u w=0.5u l=0.13u
X90 VPWR a_620_930# a_656_351# VPWR sg13_lv_pmos ad=0.104p pd=1.34u as=59f ps=0.74u w=0.2u l=0.13u
X91 Vout VGND cap_cmim l=6.99u w=6.99u
X92 a_4710_n1958# vctl VGND VGND sg13_lv_nmos ad=65.99999f pd=0.74u as=0.102p ps=1.28u w=0.3u l=0.13u
X93 a_3368_n1958# a_3429_n2395# a_2087_n2395# VGND sg13_lv_nmos ad=0.17p pd=1.68u as=0.11p ps=0.94u w=0.5u l=0.13u
X94 a_3340_351# a_2092_351# a_3434_351# VPWR sg13_lv_pmos ad=0.17p pd=1.68u as=0.11p ps=0.94u w=0.5u l=0.13u
X95 a_4709_n2525# a_620_930# VPWR VPWR sg13_lv_pmos ad=59.75f pd=0.745u as=59f ps=0.74u w=0.2u l=0.13u
X96 a_4771_n2395# a_6113_n2395# a_6052_n1958# VGND sg13_lv_nmos ad=0.11p pd=0.94u as=0.17p ps=1.68u w=0.5u l=0.13u
X97 a_656_351# a_542_269# a_750_351# VPWR sg13_lv_pmos ad=0.11p pd=0.94u as=0.1106p ps=0.945u w=0.5u l=0.13u
X98 a_2087_n2395# VGND cap_cmim l=6.99u w=6.99u
X99 VGND vctl a_620_930# VGND sg13_lv_nmos ad=0.102p pd=1.28u as=65.99999f ps=0.74u w=0.3u l=0.13u
X100 Vout a_4776_351# a_6024_351# VPWR sg13_lv_pmos ad=0.1106p pd=0.945u as=0.17p ps=1.68u w=0.5u l=0.13u
X101 a_2092_351# VGND cap_cmim l=6.99u w=6.99u
X102 a_4709_n2525# a_4771_n2395# a_3429_n2395# VPWR sg13_lv_pmos ad=0.17p pd=1.68u as=0.1106p ps=0.945u w=0.5u l=0.13u
X103 VPWR a_620_930# a_620_930# VPWR sg13_lv_pmos ad=0.104p pd=1.34u as=59.75f ps=0.745u w=0.2u l=0.13u
X104 a_4776_351# a_3434_351# a_4682_351# VPWR sg13_lv_pmos ad=0.11p pd=0.94u as=0.11p ps=0.94u w=0.5u l=0.13u
X105 a_750_351# VGND cap_cmim l=6.99u w=6.99u
X106 VGND vctl a_3368_n1958# VGND sg13_lv_nmos ad=0.102p pd=1.28u as=65.99999f ps=0.74u w=0.3u l=0.13u
X107 a_4709_n2525# a_620_930# VPWR VPWR sg13_lv_pmos ad=59f pd=0.74u as=0.104p ps=1.34u w=0.2u l=0.13u
X108 VPWR a_620_930# a_683_n2525# VPWR sg13_lv_pmos ad=0.104p pd=1.34u as=59.75f ps=0.745u w=0.2u l=0.13u
X109 a_7397_n2523# a_620_930# VPWR VPWR sg13_lv_pmos ad=59.75f pd=0.745u as=59f ps=0.74u w=0.2u l=0.13u
X110 a_683_n2525# a_745_n2395# a_542_269# VPWR sg13_lv_pmos ad=0.17p pd=1.68u as=0.1106p ps=0.945u w=0.5u l=0.13u
X111 a_4776_351# a_3434_351# a_4682_351# VPWR sg13_lv_pmos ad=0.1106p pd=0.945u as=0.17p ps=1.68u w=0.5u l=0.13u
X112 a_6052_n1958# vctl VGND VGND sg13_lv_nmos ad=65.99999f pd=0.74u as=0.102p ps=1.28u w=0.3u l=0.13u
X113 a_6113_n2395# VGND cap_cmim l=6.99u w=6.99u
X114 a_620_930# a_620_930# VPWR VPWR sg13_lv_pmos ad=59.75f pd=0.745u as=59f ps=0.74u w=0.2u l=0.13u
X115 a_2026_n1958# a_2087_n2395# a_745_n2395# VGND sg13_lv_nmos ad=0.17p pd=1.68u as=0.11p ps=0.94u w=0.5u l=0.13u
X116 a_6024_351# a_4776_351# Vout VPWR sg13_lv_pmos ad=0.11p pd=0.94u as=0.1106p ps=0.945u w=0.5u l=0.13u
X117 a_6051_n2525# a_620_930# VPWR VPWR sg13_lv_pmos ad=59.75f pd=0.745u as=59f ps=0.74u w=0.2u l=0.13u
X118 a_4710_n1958# a_4771_n2395# a_3429_n2395# VGND sg13_lv_nmos ad=0.17p pd=1.68u as=0.11p ps=0.94u w=0.5u l=0.13u
X119 a_745_n2395# VGND cap_cmim l=6.99u w=6.99u
X120 a_750_351# a_542_269# a_656_351# VPWR sg13_lv_pmos ad=0.11p pd=0.94u as=0.11p ps=0.94u w=0.5u l=0.13u
X121 a_4776_351# VGND cap_cmim l=6.99u w=6.99u
X122 VPWR a_620_930# a_1998_351# VPWR sg13_lv_pmos ad=0.104p pd=1.34u as=59f ps=0.74u w=0.2u l=0.13u
X123 a_7397_n2523# Vout a_6113_n2395# VPWR sg13_lv_pmos ad=0.11p pd=0.94u as=0.11p ps=0.94u w=0.5u l=0.13u
X124 VGND vctl a_2026_n1958# VGND sg13_lv_nmos ad=0.102p pd=1.28u as=65.99999f ps=0.74u w=0.3u l=0.13u
X125 a_1998_351# a_620_930# VPWR VPWR sg13_lv_pmos ad=59.75f pd=0.745u as=0.104p ps=1.34u w=0.2u l=0.13u
X126 a_3367_n2525# a_620_930# VPWR VPWR sg13_lv_pmos ad=59f pd=0.74u as=0.104p ps=1.34u w=0.2u l=0.13u
X127 a_2087_n2395# a_3429_n2395# a_3367_n2525# VPWR sg13_lv_pmos ad=0.11p pd=0.94u as=0.17p ps=1.68u w=0.5u l=0.13u
X128 VGND vctl a_4710_n1958# VGND sg13_lv_nmos ad=0.102p pd=1.28u as=65.99999f ps=0.74u w=0.3u l=0.13u
X129 a_3340_351# a_620_930# VPWR VPWR sg13_lv_pmos ad=59f pd=0.74u as=59f ps=0.74u w=0.2u l=0.13u
X130 a_750_351# a_542_269# a_656_351# VPWR sg13_lv_pmos ad=0.1106p pd=0.945u as=0.17p ps=1.68u w=0.5u l=0.13u
X131 a_750_351# a_542_269# a_883_n217# VGND sg13_lv_nmos ad=0.11p pd=0.94u as=0.17p ps=1.68u w=0.5u l=0.13u
X132 a_883_n217# vctl VGND VGND sg13_lv_nmos ad=65.99999f pd=0.74u as=0.102p ps=1.28u w=0.3u l=0.13u
X133 Vout a_4776_351# a_6024_351# VPWR sg13_lv_pmos ad=0.11p pd=0.94u as=0.11p ps=0.94u w=0.5u l=0.13u
X134 VPWR a_620_930# a_4682_351# VPWR sg13_lv_pmos ad=59f pd=0.74u as=59.75f ps=0.745u w=0.2u l=0.13u
X135 a_6024_351# a_620_930# VPWR VPWR sg13_lv_pmos ad=59f pd=0.74u as=59f ps=0.74u w=0.2u l=0.13u
X136 VPWR a_620_930# a_683_n2525# VPWR sg13_lv_pmos ad=59f pd=0.74u as=59f ps=0.74u w=0.2u l=0.13u
X137 a_3429_n2395# a_4771_n2395# a_4709_n2525# VPWR sg13_lv_pmos ad=0.1106p pd=0.945u as=0.11p ps=0.94u w=0.5u l=0.13u
X138 a_683_n2525# a_745_n2395# a_542_269# VPWR sg13_lv_pmos ad=0.11p pd=0.94u as=0.11p ps=0.94u w=0.5u l=0.13u
X139 a_1998_351# a_750_351# a_2092_351# VPWR sg13_lv_pmos ad=0.11p pd=0.94u as=0.1106p ps=0.945u w=0.5u l=0.13u
X140 a_6113_n2395# Vout a_7398_n1956# VGND sg13_lv_nmos ad=0.11p pd=0.94u as=0.17p ps=1.68u w=0.5u l=0.13u
X141 a_656_351# a_620_930# VPWR VPWR sg13_lv_pmos ad=59f pd=0.74u as=59f ps=0.74u w=0.2u l=0.13u
X142 VPWR a_620_930# a_7397_n2523# VPWR sg13_lv_pmos ad=0.104p pd=1.34u as=59.75f ps=0.745u w=0.2u l=0.13u
X143 VPWR a_620_930# a_2025_n2525# VPWR sg13_lv_pmos ad=59f pd=0.74u as=59f ps=0.74u w=0.2u l=0.13u
X144 VPWR a_620_930# a_1998_351# VPWR sg13_lv_pmos ad=59f pd=0.74u as=59.75f ps=0.745u w=0.2u l=0.13u
X145 a_745_n2395# a_2087_n2395# a_2026_n1958# VGND sg13_lv_nmos ad=0.11p pd=0.94u as=0.17p ps=1.68u w=0.5u l=0.13u
X146 a_3567_n217# a_2092_351# a_3434_351# VGND sg13_lv_nmos ad=0.17p pd=1.68u as=0.11p ps=0.94u w=0.5u l=0.13u
X147 VGND vctl a_3567_n217# VGND sg13_lv_nmos ad=0.102p pd=1.28u as=65.99999f ps=0.74u w=0.3u l=0.13u
X148 a_3429_n2395# a_4771_n2395# a_4709_n2525# VPWR sg13_lv_pmos ad=0.11p pd=0.94u as=0.17p ps=1.68u w=0.5u l=0.13u
C0 vctl a_4909_n217# 0.08436f
C1 a_2092_351# a_1998_351# 0.42202f
C2 a_620_930# a_6051_n2525# 0.19288f
C3 a_683_n2525# a_745_n2395# 0.10818f
C4 a_620_930# a_7397_n2523# 0.19389f
C5 VPWR a_3567_n217# 0.0108f
C6 a_2087_n2395# a_2026_n1958# 0.03943f
C7 a_2025_n2525# a_620_930# 0.18981f
C8 Vout a_6052_n1958# 0.02056f
C9 a_883_n217# a_542_269# 0.03491f
C10 VPWR Vout 0.98762f
C11 a_3429_n2395# vctl 0.04109f
C12 vctl m6_8408_n599# 0.01477f
C13 a_2087_n2395# a_2025_n2525# 0.12991f
C14 a_3429_n2395# a_620_930# 0.04637f
C15 a_7398_n1956# vctl 0.05123f
C16 vctl a_4771_n2395# 0.03129f
C17 a_3429_n2395# a_2087_n2395# 0.72984f
C18 VPWR a_1998_351# 1.37065f
C19 a_7398_n1956# a_620_930# 0.01439f
C20 VPWR a_542_269# 0.7984f
C21 a_4771_n2395# a_620_930# 0.04406f
C22 a_3434_351# a_4682_351# 0.09926f
C23 Vout a_6113_n2395# 0.81343f
C24 a_6052_n1958# a_6113_n2395# 0.03243f
C25 a_3434_351# a_4909_n217# 0.03153f
C26 VPWR a_6113_n2395# 1.36426f
C27 vctl a_4710_n1958# 0.05026f
C28 Vout a_6024_351# 0.4131f
C29 VPWR a_6024_351# 1.36969f
C30 VPWR a_4682_351# 1.35049f
C31 a_3429_n2395# a_3367_n2525# 0.12854f
C32 a_3429_n2395# a_4709_n2525# 0.45955f
C33 VPWR a_2026_n1958# 0.01457f
C34 VPWR a_6051_n2525# 1.38336f
C35 vctl a_745_n2395# 0.04038f
C36 Vout a_7397_n2523# 0.11621f
C37 VPWR a_7397_n2523# 1.38295f
C38 a_3368_n1958# vctl 0.05041f
C39 a_2225_n217# a_750_351# 0.03153f
C40 VPWR a_2025_n2525# 1.36925f
C41 a_745_n2395# a_620_930# 0.08011f
C42 a_656_351# a_750_351# 0.42803f
C43 a_4771_n2395# a_4709_n2525# 0.11922f
C44 a_745_n2395# a_684_n1958# 0.04971f
C45 a_2087_n2395# a_745_n2395# 0.35714f
C46 vctl a_750_351# 0.02282f
C47 a_683_n2525# a_620_930# 0.23019f
C48 a_3429_n2395# VPWR 1.08631f
C49 a_3368_n1958# a_2087_n2395# 0.23444f
C50 m6_8408_n599# Vout 0.01121f
C51 VPWR m6_8408_n599# 0.01344f
C52 a_750_351# a_620_930# 0.08218f
C53 a_2087_n2395# a_683_n2525# 0.01232f
C54 a_6251_n217# a_4776_351# 0.03205f
C55 a_7398_n1956# Vout 0.13041f
C56 a_4771_n2395# a_6052_n1958# 0.22936f
C57 a_4771_n2395# VPWR 0.98193f
C58 a_6113_n2395# a_6051_n2525# 0.10827f
C59 a_7397_n2523# a_6113_n2395# 0.46077f
C60 vctl a_4776_351# 0.026f
C61 a_4776_351# a_620_930# 0.04298f
C62 a_750_351# a_2092_351# 0.77984f
C63 a_6251_n217# vctl 0.08336f
C64 a_883_n217# a_750_351# 0.22378f
C65 vctl a_2225_n217# 0.07714f
C66 a_7398_n1956# a_6113_n2395# 0.21632f
C67 a_4771_n2395# a_6113_n2395# 0.58365f
C68 VPWR a_745_n2395# 0.81739f
C69 a_3368_n1958# VPWR 0.01475f
C70 a_656_351# a_620_930# 0.24146f
C71 VPWR a_683_n2525# 1.35573f
C72 vctl a_620_930# 0.09057f
C73 a_4771_n2395# a_6051_n2525# 0.46167f
C74 VPWR a_750_351# 1.05125f
C75 vctl a_684_n1958# 0.04284f
C76 a_745_n2395# a_542_269# 0.40206f
C77 vctl a_2087_n2395# 0.04184f
C78 a_4776_351# a_3434_351# 0.91818f
C79 a_684_n1958# a_620_930# 0.06371f
C80 a_2087_n2395# a_620_930# 0.05403f
C81 a_683_n2525# a_542_269# 0.45412f
C82 a_2225_n217# a_2092_351# 0.22378f
C83 a_3429_n2395# a_4771_n2395# 0.7336f
C84 a_750_351# a_1998_351# 0.09188f
C85 a_750_351# a_542_269# 0.3548f
C86 Vout a_4776_351# 0.20831f
C87 VPWR a_4776_351# 1.09569f
C88 vctl a_2092_351# 0.0248f
C89 a_3340_351# a_620_930# 0.19603f
C90 a_2026_n1958# a_745_n2395# 0.23834f
C91 a_2092_351# a_620_930# 0.04f
C92 vctl a_883_n217# 0.08086f
C93 a_3429_n2395# a_4710_n1958# 0.23035f
C94 a_620_930# a_3367_n2525# 0.19098f
C95 a_883_n217# a_620_930# 0.02036f
C96 vctl a_3434_351# 0.02497f
C97 a_620_930# a_4709_n2525# 0.18962f
C98 a_6251_n217# Vout 0.2448f
C99 a_2025_n2525# a_745_n2395# 0.42019f
C100 a_3434_351# a_620_930# 0.04103f
C101 VPWR a_2225_n217# 0.01623f
C102 VPWR a_656_351# 1.37421f
C103 a_2087_n2395# a_3367_n2525# 0.45379f
C104 vctl a_3567_n217# 0.0811f
C105 a_4771_n2395# a_4710_n1958# 0.03159f
C106 a_3429_n2395# a_3368_n1958# 0.03778f
C107 vctl Vout 0.21825f
C108 vctl a_6052_n1958# 0.04998f
C109 vctl VPWR 0.2823f
C110 a_2092_351# a_3340_351# 0.10275f
C111 Vout a_620_930# 0.16863f
C112 VPWR a_620_930# 13.1862f
C113 a_4776_351# a_6024_351# 0.1057f
C114 a_4776_351# a_4682_351# 0.42665f
C115 a_656_351# a_542_269# 0.08875f
C116 VPWR a_2087_n2395# 1.15543f
C117 a_3434_351# a_3340_351# 0.42148f
C118 a_4776_351# a_4909_n217# 0.22378f
C119 a_3434_351# a_2092_351# 0.88103f
C120 a_620_930# a_1998_351# 0.19723f
C121 a_542_269# a_620_930# 0.93638f
C122 a_3567_n217# a_2092_351# 0.03153f
C123 vctl a_6113_n2395# 0.02267f
C124 VPWR a_3340_351# 1.36686f
C125 a_684_n1958# a_542_269# 0.23665f
C126 VPWR a_2092_351# 1.29553f
C127 a_620_930# a_6113_n2395# 0.06975f
C128 m6_8408_n599# a_4776_351# 0.08511f
C129 VPWR a_3367_n2525# 1.37334f
C130 a_3567_n217# a_3434_351# 0.22378f
C131 VPWR a_4709_n2525# 1.36202f
C132 a_6024_351# a_620_930# 0.10045f
C133 vctl a_2026_n1958# 0.04894f
C134 a_4682_351# a_620_930# 0.19696f
C135 VPWR a_3434_351# 1.00449f
R0 Vout.n4 Vout.n0 30.5219
R1 Vout.n3 Vout.n1 15.6071
R2 Vout.n3 Vout.n2 15.0005
R3 Vout Vout.n4 13.4994
R4 Vout.n4 Vout.n3 9.03447
R5 vctl.n22 vctl.n0 33.8794
R6 vctl.n21 vctl.n20 33.5376
R7 vctl.n6 vctl.n4 24.4981
R8 vctl.n10 vctl.n9 24.4978
R9 vctl.n14 vctl.n13 24.4978
R10 vctl.n18 vctl.n17 24.495
R11 vctl.n6 vctl.n5 24.4894
R12 vctl.n10 vctl.n8 24.488
R13 vctl.n18 vctl.n16 24.4838
R14 vctl.n14 vctl.n12 24.4796
R15 vctl.n3 vctl.n1 24.4574
R16 vctl.n3 vctl.n2 24.4469
R17 vctl.n7 vctl.n3 10.719
R18 vctl.n19 vctl.n18 9.0005
R19 vctl.n15 vctl.n14 9.0005
R20 vctl.n11 vctl.n10 9.0005
R21 vctl.n7 vctl.n6 9.0005
R22 vctl.n21 vctl.n19 1.69764
R23 vctl.n19 vctl.n15 1.68884
R24 vctl.n15 vctl.n11 1.68004
R25 vctl.n11 vctl.n7 1.66496
R26 vctl vctl.n22 0.698214
R27 vctl.n22 vctl.n21 0.569986
R28 VGND.n94 VGND.n50 795000
R29 VGND.n92 VGND.n63 408611
R30 VGND.n84 VGND.n7 33779.7
R31 VGND.n79 VGND.n77 27000
R32 VGND.n77 VGND.n76 27000
R33 VGND.n89 VGND.n88 24089.8
R34 VGND.n91 VGND.n90 24089.8
R35 VGND.n93 VGND.n92 22334.8
R36 VGND.n87 VGND.n86 21736.5
R37 VGND.n93 VGND.n62 21565.7
R38 VGND.n84 VGND.n83 18914.1
R39 VGND.n83 VGND.n82 16059.5
R40 VGND.n85 VGND.n7 14324.5
R41 VGND.n82 VGND.n80 12933.5
R42 VGND.n169 VGND.n7 11796.7
R43 VGND.n77 VGND.n66 6755.73
R44 VGND.n77 VGND.n67 6755.73
R45 VGND.n76 VGND.n68 6755.73
R46 VGND.n79 VGND.n78 6755.73
R47 VGND.n89 VGND.n28 6068.7
R48 VGND.n90 VGND.n64 6068.7
R49 VGND.n91 VGND.n39 6068.7
R50 VGND.n88 VGND.n65 6068.7
R51 VGND.n87 VGND.n17 6068.7
R52 VGND.n86 VGND.n85 5966.17
R53 VGND.n63 VGND.n62 5388.03
R54 VGND.n75 VGND.n74 5194.39
R55 VGND.n76 VGND.n75 4867.89
R56 VGND.n80 VGND.n66 4736.52
R57 VGND.n94 VGND.n93 3958.31
R58 VGND.n64 VGND.n63 3571.26
R59 VGND.n80 VGND.n79 3511.59
R60 VGND.n75 VGND.n66 3126.84
R61 VGND.n95 VGND.n94 3045.98
R62 VGND.n85 VGND.n65 2384.11
R63 VGND.n65 VGND.n64 2380.84
R64 VGND.n82 VGND.n81 1739.46
R65 VGND.n163 VGND.n15 1155.83
R66 VGND.n148 VGND.n26 1155.83
R67 VGND.n133 VGND.n37 1155.83
R68 VGND.n118 VGND.n48 1155.83
R69 VGND.n95 VGND.n62 303.187
R70 VGND.n8 VGND.n6 295.596
R71 VGND.n162 VGND.n17 281.534
R72 VGND.n78 VGND.n23 281.534
R73 VGND.n147 VGND.n28 281.534
R74 VGND.n67 VGND.n34 281.534
R75 VGND.n132 VGND.n39 281.534
R76 VGND.n68 VGND.n45 281.534
R77 VGND.n96 VGND.n56 259.877
R78 VGND.n74 VGND.n73 258.904
R79 VGND.n117 VGND.n50 113.647
R80 VGND.n96 VGND.n95 113.186
R81 VGND.n83 VGND.n12 112.356
R82 VGND.n73 VGND.n50 108.234
R83 VGND.n56 VGND.n50 108.23
R84 VGND.n8 VGND.n5 81.1713
R85 VGND.n170 VGND.n6 76.6465
R86 VGND.n86 VGND.n84 40.634
R87 VGND.n170 VGND.n169 18.3095
R88 VGND.n90 VGND.n89 17.9646
R89 VGND.n92 VGND.n91 17.9646
R90 VGND.n88 VGND.n87 17.9646
R91 VGND.n104 VGND.n103 17.0177
R92 VGND.n161 VGND.n160 17.0005
R93 VGND.n146 VGND.n145 17.0005
R94 VGND.n131 VGND.n130 17.0005
R95 VGND.n116 VGND.n115 17.0005
R96 VGND.n110 VGND.n46 9.08291
R97 VGND.n107 VGND.n52 9.08291
R98 VGND.n125 VGND.n35 9.08291
R99 VGND.n122 VGND.n41 9.08291
R100 VGND.n140 VGND.n24 9.08291
R101 VGND.n137 VGND.n30 9.08291
R102 VGND.n155 VGND.n13 9.08291
R103 VGND.n152 VGND.n19 9.08291
R104 VGND.n97 VGND.n57 9.08291
R105 VGND.n71 VGND.n69 9.07736
R106 VGND.n3 VGND.n0 9.03039
R107 VGND VGND.n173 9.02847
R108 VGND.n109 VGND.n108 9.0005
R109 VGND.n112 VGND.n111 9.0005
R110 VGND.n124 VGND.n123 9.0005
R111 VGND.n127 VGND.n126 9.0005
R112 VGND.n139 VGND.n138 9.0005
R113 VGND.n142 VGND.n141 9.0005
R114 VGND.n154 VGND.n153 9.0005
R115 VGND.n157 VGND.n156 9.0005
R116 VGND.n102 VGND.n101 9.0005
R117 VGND.n99 VGND.n98 9.0005
R118 VGND.n100 VGND.n59 9.0005
R119 VGND.n70 VGND.n61 9.0005
R120 VGND.n113 VGND.n54 9.0005
R121 VGND.n128 VGND.n43 9.0005
R122 VGND.n143 VGND.n32 9.0005
R123 VGND.n158 VGND.n21 9.0005
R124 VGND.n160 VGND.n159 9.0005
R125 VGND.n145 VGND.n144 9.0005
R126 VGND.n130 VGND.n129 9.0005
R127 VGND.n115 VGND.n114 9.0005
R128 VGND.n2 VGND.n1 9.0005
R129 VGND.n173 VGND.n172 9.0005
R130 VGND.n81 VGND.n9 8.5005
R131 VGND.n72 VGND.n60 8.4728
R132 VGND.n104 VGND.n58 8.4706
R133 VGND.n116 VGND.n53 8.4706
R134 VGND.n131 VGND.n42 8.4706
R135 VGND.n146 VGND.n31 8.4706
R136 VGND.n161 VGND.n20 8.4706
R137 VGND.n72 VGND.n71 5.63627
R138 VGND.n119 VGND.n47 5.63396
R139 VGND.n134 VGND.n36 5.63396
R140 VGND.n149 VGND.n25 5.63396
R141 VGND.n164 VGND.n14 5.63396
R142 VGND.n119 VGND.n46 5.63382
R143 VGND.n116 VGND.n52 5.63382
R144 VGND.n134 VGND.n35 5.63382
R145 VGND.n131 VGND.n41 5.63382
R146 VGND.n149 VGND.n24 5.63382
R147 VGND.n146 VGND.n30 5.63382
R148 VGND.n164 VGND.n13 5.63382
R149 VGND.n161 VGND.n19 5.63382
R150 VGND.n104 VGND.n57 5.63382
R151 VGND.n140 VGND.n27 5.40173
R152 VGND.n97 VGND.n96 5.39607
R153 VGND.n155 VGND.n16 5.39516
R154 VGND.n125 VGND.n38 5.39516
R155 VGND.n110 VGND.n49 5.39513
R156 VGND.n74 VGND.n69 5.36707
R157 VGND.n152 VGND.n18 5.3654
R158 VGND.n137 VGND.n29 5.3654
R159 VGND.n122 VGND.n40 5.3654
R160 VGND.n107 VGND.n51 5.3654
R161 VGND.n15 VGND.n12 5.16623
R162 VGND.n163 VGND.n162 5.16623
R163 VGND.n26 VGND.n23 5.16623
R164 VGND.n148 VGND.n147 5.16623
R165 VGND.n37 VGND.n34 5.16623
R166 VGND.n133 VGND.n132 5.16623
R167 VGND.n48 VGND.n45 5.16623
R168 VGND.n118 VGND.n117 5.16623
R169 VGND VGND.n0 4.5188
R170 VGND.n78 VGND.n17 3.8748
R171 VGND.n67 VGND.n28 3.8748
R172 VGND.n68 VGND.n39 3.8748
R173 VGND.n81 VGND.n5 3.38905
R174 VGND.n172 VGND.n171 3.12829
R175 VGND.n105 VGND.n104 2.95625
R176 VGND.n165 VGND.n164 2.95625
R177 VGND.n150 VGND.n149 2.95625
R178 VGND.n135 VGND.n134 2.95625
R179 VGND.n120 VGND.n119 2.95625
R180 VGND.n161 VGND.n11 2.9562
R181 VGND.n146 VGND.n22 2.9562
R182 VGND.n131 VGND.n33 2.9562
R183 VGND.n116 VGND.n44 2.9562
R184 VGND.n10 VGND.n9 2.9539
R185 VGND.n171 VGND.n5 2.83458
R186 VGND.n163 VGND.n16 2.83383
R187 VGND.n16 VGND.n12 2.83383
R188 VGND.n148 VGND.n27 2.83383
R189 VGND.n27 VGND.n23 2.83383
R190 VGND.n133 VGND.n38 2.83383
R191 VGND.n38 VGND.n34 2.83383
R192 VGND.n118 VGND.n49 2.83383
R193 VGND.n49 VGND.n45 2.83383
R194 VGND.n162 VGND.n18 2.83383
R195 VGND.n18 VGND.n15 2.83383
R196 VGND.n147 VGND.n29 2.83383
R197 VGND.n29 VGND.n26 2.83383
R198 VGND.n132 VGND.n40 2.83383
R199 VGND.n40 VGND.n37 2.83383
R200 VGND.n117 VGND.n51 2.83383
R201 VGND.n51 VGND.n48 2.83383
R202 VGND.n164 VGND.n12 2.83383
R203 VGND.n149 VGND.n23 2.83383
R204 VGND.n134 VGND.n34 2.83383
R205 VGND.n119 VGND.n45 2.83383
R206 VGND.n119 VGND.n118 2.83383
R207 VGND.n134 VGND.n133 2.83383
R208 VGND.n149 VGND.n148 2.83383
R209 VGND.n164 VGND.n163 2.83383
R210 VGND.n161 VGND.n15 2.83383
R211 VGND.n162 VGND.n161 2.83383
R212 VGND.n146 VGND.n26 2.83383
R213 VGND.n147 VGND.n146 2.83383
R214 VGND.n131 VGND.n37 2.83383
R215 VGND.n132 VGND.n131 2.83383
R216 VGND.n116 VGND.n48 2.83383
R217 VGND.n117 VGND.n116 2.83383
R218 VGND.n171 VGND.n170 2.83383
R219 VGND.n171 VGND.n4 2.80958
R220 VGND.n167 VGND.n9 2.73145
R221 VGND.n168 VGND.n167 2.6007
R222 VGND.n72 VGND.n55 2.48001
R223 VGND.n4 VGND.n3 0.962312
R224 VGND.n169 VGND.n168 0.744345
R225 VGND.n114 VGND.n113 0.3701
R226 VGND.n129 VGND.n128 0.3701
R227 VGND.n144 VGND.n143 0.3701
R228 VGND.n159 VGND.n158 0.3701
R229 VGND.n101 VGND.n100 0.3701
R230 VGND.n172 VGND.n2 0.3555
R231 VGND.n3 VGND.n2 0.353
R232 VGND.n166 VGND.n10 0.325527
R233 VGND.n21 VGND.n11 0.323287
R234 VGND.n32 VGND.n22 0.323287
R235 VGND.n43 VGND.n33 0.323287
R236 VGND.n54 VGND.n44 0.323287
R237 VGND.n103 VGND.n55 0.262968
R238 VGND.n167 VGND.n166 0.223793
R239 VGND.n10 VGND.n4 0.195252
R240 VGND.n109 VGND.n107 0.192746
R241 VGND.n112 VGND.n110 0.192746
R242 VGND.n124 VGND.n122 0.192746
R243 VGND.n127 VGND.n125 0.192746
R244 VGND.n139 VGND.n137 0.192746
R245 VGND.n142 VGND.n140 0.192746
R246 VGND.n154 VGND.n152 0.192746
R247 VGND.n157 VGND.n155 0.192746
R248 VGND.n69 VGND.n61 0.192746
R249 VGND.n99 VGND.n97 0.192746
R250 VGND.n114 VGND.n109 0.191392
R251 VGND.n113 VGND.n112 0.191392
R252 VGND.n129 VGND.n124 0.191392
R253 VGND.n128 VGND.n127 0.191392
R254 VGND.n144 VGND.n139 0.191392
R255 VGND.n143 VGND.n142 0.191392
R256 VGND.n159 VGND.n154 0.191392
R257 VGND.n158 VGND.n157 0.191392
R258 VGND.n101 VGND.n61 0.191392
R259 VGND.n100 VGND.n99 0.191392
R260 VGND.n108 VGND.n52 0.163122
R261 VGND.n123 VGND.n41 0.163122
R262 VGND.n138 VGND.n30 0.163122
R263 VGND.n153 VGND.n19 0.163122
R264 VGND.n98 VGND.n57 0.163122
R265 VGND.n156 VGND.n13 0.163122
R266 VGND.n141 VGND.n24 0.163122
R267 VGND.n126 VGND.n35 0.163122
R268 VGND.n111 VGND.n46 0.163122
R269 VGND.n166 VGND.n165 0.161915
R270 VGND.n121 VGND.n120 0.158669
R271 VGND.n136 VGND.n135 0.158669
R272 VGND.n151 VGND.n150 0.158669
R273 VGND.n106 VGND.n105 0.158669
R274 VGND.n111 VGND.n47 0.154735
R275 VGND.n126 VGND.n36 0.154735
R276 VGND.n141 VGND.n25 0.154735
R277 VGND.n156 VGND.n14 0.154735
R278 VGND.n71 VGND.n70 0.15113
R279 VGND.n108 VGND.n53 0.123672
R280 VGND.n123 VGND.n42 0.123672
R281 VGND.n138 VGND.n31 0.123672
R282 VGND.n153 VGND.n20 0.123672
R283 VGND.n98 VGND.n58 0.123672
R284 VGND.n59 VGND.n58 0.120235
R285 VGND.n70 VGND.n60 0.114798
R286 VGND.n102 VGND.n60 0.111609
R287 VGND.n106 VGND.n53 0.0927349
R288 VGND.n121 VGND.n42 0.0927349
R289 VGND.n136 VGND.n31 0.0927349
R290 VGND.n151 VGND.n20 0.0927349
R291 VGND.n54 VGND.n47 0.06234
R292 VGND.n43 VGND.n36 0.06234
R293 VGND.n32 VGND.n25 0.06234
R294 VGND.n21 VGND.n14 0.06234
R295 VGND.n173 VGND.n1 0.0597227
R296 VGND.n105 VGND.n55 0.0487297
R297 VGND.n103 VGND.n59 0.04175
R298 VGND.n103 VGND.n102 0.0403551
R299 VGND.n1 VGND.n0 0.0302293
R300 VGND.n168 VGND.n6 0.00732966
R301 VGND.n165 VGND.n11 0.00274058
R302 VGND.n150 VGND.n22 0.00274058
R303 VGND.n135 VGND.n33 0.00274058
R304 VGND.n120 VGND.n44 0.00274058
R305 VGND.n160 VGND.n21 0.00194262
R306 VGND.n145 VGND.n32 0.00194262
R307 VGND.n130 VGND.n43 0.00194262
R308 VGND.n115 VGND.n54 0.00194262
R309 VGND.n9 VGND.n8 0.00153443
R310 VGND.n73 VGND.n72 0.00143734
R311 VGND.n104 VGND.n56 0.00111193
R312 VGND.n160 VGND.n151 0.000860656
R313 VGND.n145 VGND.n136 0.000860656
R314 VGND.n130 VGND.n121 0.000860656
R315 VGND.n115 VGND.n106 0.000860656
C136 vctl VGND 11.2448f
C137 Vout VGND 7.04733f
C138 VPWR VGND 11.0209f
C139 m6_8408_n599# VGND 1.85457f
C140 a_7397_n2523# VGND 0.05072f $ **FLOATING
C141 a_6051_n2525# VGND 0.04654f $ **FLOATING
C142 a_4709_n2525# VGND 0.0474f $ **FLOATING
C143 a_3367_n2525# VGND 0.04814f $ **FLOATING
C144 a_2025_n2525# VGND 0.04567f $ **FLOATING
C145 a_683_n2525# VGND 0.07408f $ **FLOATING
C146 a_6113_n2395# VGND 4.52843f $ **FLOATING
C147 a_4771_n2395# VGND 4.66244f $ **FLOATING
C148 a_3429_n2395# VGND 4.71205f $ **FLOATING
C149 a_2087_n2395# VGND 5.15226f $ **FLOATING
C150 a_745_n2395# VGND 5.27135f $ **FLOATING
C151 a_7398_n1956# VGND 0.75149f $ **FLOATING
C152 a_6052_n1958# VGND 0.8045f $ **FLOATING
C153 a_4710_n1958# VGND 0.81785f $ **FLOATING
C154 a_3368_n1958# VGND 0.82955f $ **FLOATING
C155 a_2026_n1958# VGND 0.82862f $ **FLOATING
C156 a_684_n1958# VGND 0.83893f $ **FLOATING
C157 a_6251_n217# VGND 0.65187f $ **FLOATING
C158 a_4909_n217# VGND 0.67139f $ **FLOATING
C159 a_3567_n217# VGND 0.6715f $ **FLOATING
C160 a_2225_n217# VGND 0.67644f $ **FLOATING
C161 a_883_n217# VGND 0.68389f $ **FLOATING
C162 a_4776_351# VGND 5.0221f $ **FLOATING
C163 a_3434_351# VGND 4.4055f $ **FLOATING
C164 a_2092_351# VGND 4.40424f $ **FLOATING
C165 a_750_351# VGND 4.67142f $ **FLOATING
C166 a_542_269# VGND 6.17341f $ **FLOATING
C167 a_6024_351# VGND 0.05888f $ **FLOATING
C168 a_4682_351# VGND 0.03844f $ **FLOATING
C169 a_3340_351# VGND 0.04051f $ **FLOATING
C170 a_1998_351# VGND 0.04084f $ **FLOATING
C171 a_656_351# VGND 0.05472f $ **FLOATING
C172 a_620_930# VGND 5.66202f $ **FLOATING
.ends
