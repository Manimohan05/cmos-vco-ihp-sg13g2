** sch_path: /foss/designs/iic-osic-tools/cmos-vco-ihp-sg13g2/Combined_Design/design_data/xschem/vco_wob_tb.sch
**.subckt vco_wob_tb Vout
*.opin Vout
VPWR net1 GND 1.2
vctl net2 GND 1
x1 net1 GND net2 Vout vco_wob
**** begin user architecture code
 .lib cornerMOSlv.lib mos_tt
.lib /foss/pdks/ihp-sg13g2/libs.tech/ngspice/models/cornerCAP.lib cap_typ_stat



.temp 27
.control
save all
.options maxstep=10n reltol=1e-3 abstol=1e-6
tran 50p 1u
plot v(Vout) xlimit 500n 1u
fft v(Vout)
plot db(mag(fft_v(vout))) xlimit 1Meg 100Meg
wrdata fft_output_Vcon1.txt db(mag(fft_v(vout)))
op
write vco_wob_tb.raw
.endc



**** end user architecture code
**.ends

* expanding   symbol:  vco_wob.sym # of pins=4
** sym_path: /foss/designs/iic-osic-tools/cmos-vco-ihp-sg13g2/Combined_Design/design_data/xschem/vco_wob.sym
** sch_path: /foss/designs/iic-osic-tools/cmos-vco-ihp-sg13g2/Combined_Design/design_data/xschem/vco_wob.sch
.subckt vco_wob VPWR VGND vctl Vout
*.iopin VPWR
*.iopin VGND
*.ipin vctl
*.opin Vout
XM21 mirror_pg mirror_pg VPWR VPWR sg13_lv_pmos w=0.8u l=0.13u ng=1 m=1
XM22 net1 mirror_pg VPWR VPWR sg13_lv_pmos w=0.8u l=0.13u ng=1 m=1
XM23 net2 mirror_pg VPWR VPWR sg13_lv_pmos w=0.8u l=0.13u ng=1 m=1
XM24 net3 mirror_pg VPWR VPWR sg13_lv_pmos w=0.8u l=0.13u ng=1 m=1
XM25 mirror_pg vctl VGND VGND sg13_lv_nmos w=0.6u l=0.13u ng=1 m=1
XM26 net9 vctl VGND VGND sg13_lv_nmos w=0.6u l=0.13u ng=1 m=1
XM28 net7 vctl VGND VGND sg13_lv_nmos w=0.6u l=0.13u ng=1 m=1
XM29 net13 mirror_pg VPWR VPWR sg13_lv_pmos w=0.8u l=0.13u ng=1 m=1
XM30 net12 mirror_pg VPWR VPWR sg13_lv_pmos w=0.8u l=0.13u ng=1 m=1
XM31 net10 vctl VGND VGND sg13_lv_nmos w=0.6u l=0.13u ng=1 m=1
XM32 net11 vctl VGND VGND sg13_lv_nmos w=0.6u l=0.13u ng=1 m=1
XM33 net15 mirror_pg VPWR VPWR sg13_lv_pmos w=0.8u l=0.13u ng=1 m=1
XM34 net16 mirror_pg VPWR VPWR sg13_lv_pmos w=0.8u l=0.13u ng=1 m=1
XM35 net20 vctl VGND VGND sg13_lv_nmos w=0.6u l=0.13u ng=1 m=1
XM36 net19 vctl VGND VGND sg13_lv_nmos w=0.6u l=0.13u ng=1 m=1
XM37 net24 mirror_pg VPWR VPWR sg13_lv_pmos w=0.8u l=0.13u ng=1 m=1
XM38 net23 mirror_pg VPWR VPWR sg13_lv_pmos w=0.8u l=0.13u ng=1 m=1
XM39 net21 vctl VGND VGND sg13_lv_nmos w=0.6u l=0.13u ng=1 m=1
XM40 net22 vctl VGND VGND sg13_lv_nmos w=0.6u l=0.13u ng=1 m=1
XM41 net31 mirror_pg VPWR VPWR sg13_lv_pmos w=0.8u l=0.13u ng=1 m=1
XM42 net30 mirror_pg VPWR VPWR sg13_lv_pmos w=0.8u l=0.13u ng=1 m=1
XM43 net28 vctl VGND VGND sg13_lv_nmos w=0.6u l=0.13u ng=1 m=1
XM44 net29 vctl VGND VGND sg13_lv_nmos w=0.6u l=0.13u ng=1 m=1
XM1 net8 vctl VGND VGND sg13_lv_nmos w=0.6u l=0.13u ng=1 m=1
XC12 net4 VGND cap_cmim w=6.99e-6 l=6.99e-6 m=1
XC1 net5 VGND cap_cmim w=6.99e-6 l=6.99e-6 m=1
XC2 net6 VGND cap_cmim w=6.99e-6 l=6.99e-6 m=1
XC3 net14 VGND cap_cmim w=6.99e-6 l=6.99e-6 m=1
XC4 net26 VGND cap_cmim w=6.99e-6 l=6.99e-6 m=1
XC5 net17 VGND cap_cmim w=6.99e-6 l=6.99e-6 m=1
XC6 net18 VGND cap_cmim w=6.99e-6 l=6.99e-6 m=1
XC7 net25 VGND cap_cmim w=6.99e-6 l=6.99e-6 m=1
XC8 net27 VGND cap_cmim w=6.99e-6 l=6.99e-6 m=1
XC9 net32 VGND cap_cmim w=6.99e-6 l=6.99e-6 m=1
XC10 Vout VGND cap_cmim w=6.99e-6 l=6.99e-6 m=1
x1 net1 VPWR Vout net4 VGND net9 vco_inverter
x2 net2 VPWR net4 net5 VGND net8 vco_inverter
x3 net3 VPWR net5 net6 VGND net7 vco_inverter
x4 net13 VPWR net6 net14 VGND net10 vco_inverter
x5 net12 VPWR net14 net26 VGND net11 vco_inverter
x6 net15 VPWR net26 net17 VGND net20 vco_inverter
x7 net16 VPWR net17 net18 VGND net19 vco_inverter
x8 net24 VPWR net18 net25 VGND net21 vco_inverter
x9 net23 VPWR net25 net27 VGND net22 vco_inverter
x10 net31 VPWR net27 net32 VGND net28 vco_inverter
x11 net30 VPWR net32 Vout VGND net29 vco_inverter
.ends


* expanding   symbol:  vco_inverter.sym # of pins=6
** sym_path: /foss/designs/iic-osic-tools/cmos-vco-ihp-sg13g2/Combined_Design/design_data/xschem/vco_inverter.sym
** sch_path: /foss/designs/iic-osic-tools/cmos-vco-ihp-sg13g2/Combined_Design/design_data/xschem/vco_inverter.sch
.subckt vco_inverter VPWR VPB A Y VNB VGND
*.iopin VPWR
*.iopin VGND
*.ipin A
*.opin Y
*.iopin VPB
*.iopin VNB
XM2 Y A VPWR VPB sg13_lv_pmos w=2u l=0.13u ng=1 m=1
XM1 Y A VGND VNB sg13_lv_nmos w=1u l=0.13u ng=1 m=1
.ends

.GLOBAL GND
.end
