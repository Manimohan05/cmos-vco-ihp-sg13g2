** sch_path: /foss/designs/iic-osic-tools/cmos-vco-ihp-sg13g2/design_data/xschem/vco_pex_tb.sch
**.subckt vco_pex_tb Vout
*.opin Vout
VPWR net1 GND 1.2
vctl net2 GND 1
x1 net1 GND net2 Vout vco
**** begin user architecture code
 .lib cornerMOSlv.lib mos_tt
.lib /foss/pdks/ihp-sg13g2/libs.tech/ngspice/models/cornerCAP.lib cap_typ_stat



.include /foss/designs/iic-osic-tools/cmos-vco-ihp-sg13g2/design_data/pex/vco__vco/magic_RC/vco.pex.spice
.param temp=27
.control
save all
.options maxstep=10n reltol=1e-3 abstol=1e-6
save v(Vout)
tran 100p 1u
write vco_pex.raw
plot v(Vout) xlimit 500n 1u
fft v(Vout)
let vmag = db(mag(v(Vout)))
plot vmag xlabel 'Frequency (Hz)' xlimit 1Meg 100Meg
wrdata fft_output(Vcon=1).txt vmag
.endc


**** end user architecture code
**.ends
.GLOBAL GND
.end
